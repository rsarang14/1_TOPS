module twiddle_rom_512 (
    input [7:0] addr, 
    output reg signed [15:0] wr, 
    output reg signed [15:0] wi
);
    // Roll Number: EC23I2015 - FFT Twiddle ROM (512-pt, Q15)
    always @(*) begin
        case(addr)
            8'h00: begin wr = 16'h7FFF; wi = 16'h0000; end
            8'h01: begin wr = 16'h7FFD; wi = 16'hFE6E; end
            8'h02: begin wr = 16'h7FF5; wi = 16'hFCDC; end
            8'h03: begin wr = 16'h7FE9; wi = 16'hFB4A; end
            8'h04: begin wr = 16'h7FD8; wi = 16'hF9B8; end
            8'h05: begin wr = 16'h7FC1; wi = 16'hF827; end
            8'h06: begin wr = 16'h7FA6; wi = 16'hF696; end
            8'h07: begin wr = 16'h7F86; wi = 16'hF505; end
            8'h08: begin wr = 16'h7F61; wi = 16'hF374; end
            8'h09: begin wr = 16'h7F37; wi = 16'hF1E4; end
            8'h0A: begin wr = 16'h7F09; wi = 16'hF055; end
            8'h0B: begin wr = 16'h7ED5; wi = 16'hEEC6; end
            8'h0C: begin wr = 16'h7E9C; wi = 16'hED38; end
            8'h0D: begin wr = 16'h7E5F; wi = 16'hEBAB; end
            8'h0E: begin wr = 16'h7E1C; wi = 16'hEA1E; end
            8'h0F: begin wr = 16'h7DD5; wi = 16'hE892; end
            8'h10: begin wr = 16'h7D8A; wi = 16'hE707; end
            8'h11: begin wr = 16'h7D39; wi = 16'hE57D; end
            8'h12: begin wr = 16'h7CE4; wi = 16'hE3F4; end
            8'h13: begin wr = 16'h7C89; wi = 16'hE26C; end
            8'h14: begin wr = 16'h7C2A; wi = 16'hE0E5; end
            8'h15: begin wr = 16'h7BC5; wi = 16'hDF60; end
            8'h16: begin wr = 16'h7B5D; wi = 16'hDDDC; end
            8'h17: begin wr = 16'h7AF0; wi = 16'hDC59; end
            8'h18: begin wr = 16'h7A7D; wi = 16'hDAD7; end
            8'h19: begin wr = 16'h7A06; wi = 16'hD957; end
            8'h1A: begin wr = 16'h798A; wi = 16'hD7D8; end
            8'h1B: begin wr = 16'h790A; wi = 16'hD65B; end
            8'h1C: begin wr = 16'h7884; wi = 16'hD4DF; end
            8'h1D: begin wr = 16'h77FA; wi = 16'hD365; end
            8'h1E: begin wr = 16'h776C; wi = 16'hD1EC; end
            8'h1F: begin wr = 16'h76DA; wi = 16'hD075; end
            8'h20: begin wr = 16'h7641; wi = 16'hCEFF; end
            8'h21: begin wr = 16'h75A5; wi = 16'hCD8C; end
            8'h22: begin wr = 16'h7504; wi = 16'hCC1B; end
            8'h23: begin wr = 16'h7460; wi = 16'hCAAB; end
            8'h24: begin wr = 16'h73B6; wi = 16'hC93D; end
            8'h25: begin wr = 16'h7308; wi = 16'hC7D1; end
            8'h26: begin wr = 16'h7255; wi = 16'hC667; end
            8'h27: begin wr = 16'h719E; wi = 16'hC4FF; end
            8'h28: begin wr = 16'h70E3; wi = 16'hC399; end
            8'h29: begin wr = 16'h7023; wi = 16'hC235; end
            8'h2A: begin wr = 16'h6F5F; wi = 16'hC0D4; end
            8'h2B: begin wr = 16'h6E97; wi = 16'hBF75; end
            8'h2C: begin wr = 16'h6DCA; wi = 16'hBE18; end
            8'h2D: begin wr = 16'h6CFA; wi = 16'hBCBD; end
            8'h2E: begin wr = 16'h6C24; wi = 16'hBB64; end
            8'h2F: begin wr = 16'h6B4A; wi = 16'hBA0E; end
            8'h30: begin wr = 16'h6A6D; wi = 16'hB8BA; end
            8'h31: begin wr = 16'h698C; wi = 16'hB769; end
            8'h32: begin wr = 16'h68A7; wi = 16'hB61A; end
            8'h33: begin wr = 16'h67BE; wi = 16'hB4CD; end
            8'h34: begin wr = 16'h66D1; wi = 16'hB383; end
            8'h35: begin wr = 16'h65E0; wi = 16'hB23B; end
            8'h36: begin wr = 16'h64EB; wi = 16'hB0F5; end
            8'h37: begin wr = 16'h63F3; wi = 16'hAFB3; end
            8'h38: begin wr = 16'h62F7; wi = 16'hAE73; end
            8'h39: begin wr = 16'h61F7; wi = 16'hAD35; end
            8'h3A: begin wr = 16'h60F3; wi = 16'hABF9; end
            8'h3B: begin wr = 16'h5FEB; wi = 16'hAABF; end
            8'h3C: begin wr = 16'h5EDF; wi = 16'hA988; end
            8'h3D: begin wr = 16'h5DCF; wi = 16'hA854; end
            8'h3E: begin wr = 16'h5CBB; wi = 16'hA722; end
            8'h3F: begin wr = 16'h5BA3; wi = 16'hA5F4; end
            8'h40: begin wr = 16'h5A82; wi = 16'hA57E; end
            8'h41: begin wr = 16'h595E; wi = 16'hA45D; end
            8'h42: begin wr = 16'h5836; wi = 16'hA33F; end
            8'h43: begin wr = 16'h570A; wi = 16'hA224; end
            8'h44: begin wr = 16'h55DB; wi = 16'hA111; end
            8'h45: begin wr = 16'h54A7; wi = 16'hA001; end
            8'h46: begin wr = 16'h5370; wi = 16'h9EF5; end
            8'h47: begin wr = 16'h5235; wi = 16'h9DEC; end
            8'h48: begin wr = 16'h50F5; wi = 16'h9CE7; end
            8'h49: begin wr = 16'h4FB3; wi = 16'h9BE5; end
            8'h4A: begin wr = 16'h4E6D; wi = 16'h9AE8; end
            8'h4B: begin wr = 16'h4D23; wi = 16'h99EE; end
            8'h4C: begin wr = 16'h4BD4; wi = 16'h98F9; end
            8'h4D: begin wr = 16'h4A82; wi = 16'h9807; end
            8'h4E: begin wr = 16'h492C; wi = 16'h971A; end
            8'h4F: begin wr = 16'h47D3; wi = 16'h9631; end
            8'h50: begin wr = 16'h4677; wi = 16'h954D; end
            8'h51: begin wr = 16'h4517; wi = 16'h946D; end
            8'h52: begin wr = 16'h43B5; wi = 16'h9391; end
            8'h53: begin wr = 16'h424E; wi = 16'h92B9; end
            8'h54: begin wr = 16'h40E5; wi = 16'h91E6; end
            8'h55: begin wr = 16'h3F78; wi = 16'h9118; end
            8'h56: begin wr = 16'h3E0A; wi = 16'h904D; end
            8'h57: begin wr = 16'h3C99; wi = 16'h8F88; end
            8'h58: begin wr = 16'h3B25; wi = 16'h8EC8; end
            8'h59: begin wr = 16'h39AF; wi = 16'h8E0D; end
            8'h5A: begin wr = 16'h3736; wi = 16'h8D56; end
            8'h5B: begin wr = 16'h35BA; wi = 16'h8CA5; end
            8'h5C: begin wr = 16'h343C; wi = 16'h8BF9; end
            8'h5D: begin wr = 16'h32BC; wi = 16'h8B51; end
            8'h5E: begin wr = 16'h3139; wi = 16'h8AAE; end
            8'h5F: begin wr = 16'h2FB4; wi = 16'h8A11; end
            8'h60: begin wr = 16'h2E2D; wi = 16'h8979; end
            8'h61: begin wr = 16'h2CA4; wi = 16'h88E6; end
            8'h62: begin wr = 16'h2B19; wi = 16'h885A; end
            8'h63: begin wr = 16'h298C; wi = 16'h87D4; end
            8'h64: begin wr = 16'h27FD; wi = 16'h8754; end
            8'h65: begin wr = 16'h266C; wi = 16'h86D9; end
            8'h66: begin wr = 16'h24DA; wi = 16'h8664; end
            8'h67: begin wr = 16'h2346; wi = 16'h85F5; end
            8'h68: begin wr = 16'h21B0; wi = 16'h858E; end
            8'h69: begin wr = 16'h2019; wi = 16'h852E; end
            8'h6A: begin wr = 16'h1E80; wi = 16'h84D4; end
            8'h6B: begin wr = 16'h1CE6; wi = 16'h8480; end
            8'h6C: begin wr = 16'h1B4A; wi = 16'h8433; end
            8'h6D: begin wr = 16'h19AD; wi = 16'h83EE; end
            8'h6E: begin wr = 16'h1810; wi = 16'h83B0; end
            8'h6F: begin wr = 16'h1671; wi = 16'h827C; end
            8'h70: begin wr = 16'h14D2; wi = 16'h8251; end
            8'h71: begin wr = 16'h1331; wi = 16'h822D; end
            8'h72: begin wr = 16'h1191; wi = 16'h8211; end
            8'h73: begin wr = 16'h0FEE; wi = 16'h81FA; end
            8'h74: begin wr = 16'h0E4C; wi = 16'h81EA; end
            8'h75: begin wr = 16'h0CA9; wi = 16'h81DF; end
            8'h76: begin wr = 16'h0B06; wi = 16'h81DA; end
            8'h77: begin wr = 16'h0961; wi = 16'h81DC; end
            8'h78: begin wr = 16'h07BD; wi = 16'h81E3; end
            8'h79: begin wr = 16'h0618; wi = 16'h81F1; end
            8'h7A: begin wr = 16'h0473; wi = 16'h8205; end
            8'h7B: begin wr = 16'h02CE; wi = 16'h821F; end
            8'h7C: begin wr = 16'h0129; wi = 16'h823F; end
            8'h7D: begin wr = 16'hFF83; wi = 16'h8264; end
            8'h7E: begin wr = 16'hFDDE; wi = 16'h828F; end
            8'h7F: begin wr = 16'hFC39; wi = 16'h82C0; end
            8'h80: begin wr = 16'h0000; wi = 16'h8000; end
            8'h81: begin wr = 16'hE98F; wi = 16'h82C0; end
            8'h82: begin wr = 16'hF222; wi = 16'h828F; end
            8'h83: begin wr = 16'hF07D; wi = 16'h8264; end
            8'h84: begin wr = 16'hEED7; wi = 16'h823F; end
            8'h85: begin wr = 16'hED32; wi = 16'h821F; end
            8'h86: begin wr = 16'hEB8D; wi = 16'h8205; end
            8'h87: begin wr = 16'hE9E8; wi = 16'h81F1; end
            8'h88: begin wr = 16'hE843; wi = 16'h81E3; end
            8'h89: begin wr = 16'hE69F; wi = 16'h81DC; end
            8'h8A: begin wr = 16'hE4FA; wi = 16'h81DA; end
            8'h8B: begin wr = 16'hE357; wi = 16'h81DF; end
            8'h8C: begin wr = 16'hE1B4; wi = 16'h81EA; end
            8'h8D: begin wr = 16'hE012; wi = 16'h81FA; end
            8'h8E: begin wr = 16'hDE6F; wi = 16'h8211; end
            8'h8F: begin wr = 16'hDCCF; wi = 16'h822D; end
            8'h90: begin wr = 16'hDB2E; wi = 16'h8251; end
            8'h91: begin wr = 16'hD98F; wi = 16'h827C; end
            8'h92: begin wr = 16'hD7F0; wi = 16'h83B0; end
            8'h93: begin wr = 16'hD653; wi = 16'h83EE; end
            8'h94: begin wr = 16'hD4B6; wi = 16'h8433; end
            8'h95: begin wr = 16'hD31A; wi = 16'h8480; end
            8'h96: begin wr = 16'hD180; wi = 16'h84D4; end
            8'h97: begin wr = 16'hCFE7; wi = 16'h852E; end
            8'h98: begin wr = 16'hCE50; wi = 16'h858E; end
            8'h99: begin wr = 16'hCCBA; wi = 16'h85F5; end
            8'h9A: begin wr = 16'hCB26; wi = 16'h8664; end
            8'h9B: begin wr = 16'hC994; wi = 16'h86D9; end
            8'h9C: begin wr = 16'hC803; wi = 16'h8754; end
            8'h9D: begin wr = 16'hC674; wi = 16'h87D4; end
            8'h9E: begin wr = 16'hC4E7; wi = 16'h885A; end
            8'h9F: begin wr = 16'hC35C; wi = 16'h88E6; end
            8'hA0: begin wr = 16'hC1D3; wi = 16'h8979; end
            8'hA1: begin wr = 16'hC04C; wi = 16'h8A11; end
            8'hA2: begin wr = 16'hBEC7; wi = 16'h8AAE; end
            8'hA3: begin wr = 16'hBD44; wi = 16'h8B51; end
            8'hA4: begin wr = 16'hBBC4; wi = 16'h8BF9; end
            8'hA5: begin wr = 16'hBA46; wi = 16'h8CA5; end
            8'hA6: begin wr = 16'hB8CA; wi = 16'h8D56; end
            8'hA7: begin wr = 16'hB751; wi = 16'h8E0D; end
            8'hA8: begin wr = 16'hB5DB; wi = 16'h8EC8; end
            8'hA9: begin wr = 16'hB467; wi = 16'h8F88; end
            8'hAA: begin wr = 16'hB2F6; wi = 16'h904D; end
            8'hAB: begin wr = 16'hB188; wi = 16'h9118; end
            8'hAC: begin wr = 16'hB01B; wi = 16'h91E6; end
            8'hAD: begin wr = 16'hAEB2; wi = 16'h92B9; end
            8'hAE: begin wr = 16'hAD4B; wi = 16'h9391; end
            8'hAF: begin wr = 16'hABE9; wi = 16'h946D; end
            8'hB0: begin wr = 16'hAA89; wi = 16'h954D; end
            8'hB1: begin wr = 16'hA92D; wi = 16'h9631; end
            8'hB2: begin wr = 16'hA7D4; wi = 16'h971A; end
            8'hB3: begin wr = 16'hA67E; wi = 16'h9807; end
            8'hB4: begin wr = 16'hA52C; wi = 16'h98F9; end
            8'hB5: begin wr = 16'hA3DD; wi = 16'h99EE; end
            8'hB6: begin wr = 16'hA293; wi = 16'h9AE8; end
            8'hB7: begin wr = 16'hA14D; wi = 16'h9BE5; end
            8'hB8: begin wr = 16'hA00B; wi = 16'h9CE7; end
            8'hB9: begin wr = 16'h9ECA; wi = 16'h9DEC; end
            8'hBA: begin wr = 16'h9D90; wi = 16'h9EF5; end
            8'hBB: begin wr = 16'h9C59; wi = 16'hA001; end
            8'hBC: begin wr = 16'h9B25; wi = 16'hA111; end
            8'hBD: begin wr = 16'h99F6; wi = 16'hA224; end
            8'hBE: begin wr = 16'h98CA; wi = 16'hA33F; end
            8'hBF: begin wr = 16'h97A2; wi = 16'hA45D; end
            8'hC0: begin wr = 16'h967E; wi = 16'hA57E; end
            8'hC1: begin wr = 16'h955D; wi = 16'hA5F4; end
            8'hC2: begin wr = 16'h9445; wi = 16'hA722; end
            8'hC3: begin wr = 16'h9331; wi = 16'hA854; end
            8'hC4: begin wr = 16'h9221; wi = 16'hA988; end
            8'hC5: begin wr = 16'h9115; wi = 16'hAABF; end
            8'hC6: begin wr = 16'h900D; wi = 16'hABF9; end
            8'hC7: begin wr = 16'h8F09; wi = 16'hAD35; end
            8'hC8: begin wr = 16'h8E09; wi = 16'hAE73; end
            8'hC9: begin wr = 16'h8D0D; wi = 16'hAFB3; end
            8'hCA: begin wr = 16'h8C15; wi = 16'hB0F5; end
            8'hCB: begin wr = 16'h8B20; wi = 16'hB23B; end
            8'hCC: begin wr = 16'h8A2F; wi = 16'hB383; end
            8'hCD: begin wr = 16'h8942; wi = 16'hB4CD; end
            8'hCE: begin wr = 16'h8859; wi = 16'hB61A; end
            8'hCF: begin wr = 16'h8774; wi = 16'hB769; end
            8'hD0: begin wr = 16'h8693; wi = 16'hB8BA; end
            8'hD1: begin wr = 16'h85B6; wi = 16'hBA0E; end
            8'hD2: begin wr = 16'h84DC; wi = 16'hBB64; end
            8'hD3: begin wr = 16'h8406; wi = 16'hBCBD; end
            8'hD4: begin wr = 16'h8336; wi = 16'hBE18; end
            8'hD5: begin wr = 16'h8269; wi = 16'hBF75; end
            8'hD6: begin wr = 16'h81A1; wi = 16'hC0D4; end
            8'hD7: begin wr = 16'h80DD; wi = 16'hC235; end
            8'hD8: begin wr = 16'h801D; wi = 16'hC399; end
            8'hD9: begin wr = 16'h7F62; wi = 16'hC4FF; end
            8'hDA: begin wr = 16'h7EAB; wi = 16'hC667; end
            8'hDB: begin wr = 16'h7DF8; wi = 16'hC7D1; end
            8'hDC: begin wr = 16'h7D4A; wi = 16'hC93D; end
            8'hDD: begin wr = 16'h7CA0; wi = 16'hCAAB; end
            8'hDE: begin wr = 16'h7BFC; wi = 16'hCC1B; end
            8'hDF: begin wr = 16'h7B5B; wi = 16'hCD8C; end
            8'hE0: begin wr = 16'h7ABF; wi = 16'hCEFF; end
            8'hE1: begin wr = 16'h7926; wi = 16'hD075; end
            8'hE2: begin wr = 16'h7894; wi = 16'hD1EC; end
            8'hE3: begin wr = 16'h7806; wi = 16'hD365; end
            8'hE4: begin wr = 16'h777C; wi = 16'hD4DF; end
            8'hE5: begin wr = 16'h76F6; wi = 16'hD65B; end
            8'hE6: begin wr = 16'h7676; wi = 16'hD7D8; end
            8'hE7: begin wr = 16'h75FA; wi = 16'hD957; end
            8'hE8: begin wr = 16'h7583; wi = 16'hDAD7; end
            8'hE9: begin wr = 16'h7510; wi = 16'hDC59; end
            8'hEA: begin wr = 16'h74A3; wi = 16'hDDDC; end
            8'hEB: begin wr = 16'h743B; wi = 16'hDF60; end
            8'hEC: begin wr = 16'h73D6; wi = 16'hE0E5; end
            8'hED: begin wr = 16'h7377; wi = 16'hE26C; end
            8'hEE: begin wr = 16'h731C; wi = 16'hE3F4; end
            8'hEF: begin wr = 16'h72C7; wi = 16'hE57D; end
            8'hF0: begin wr = 16'h7276; wi = 16'hE707; end
            8'hF1: begin wr = 16'h722B; wi = 16'hE892; end
            8'hF2: begin wr = 16'h71E4; wi = 16'hEA1E; end
            8'hF3: begin wr = 16'h71A1; wi = 16'hEBAB; end
            8'hF4: begin wr = 16'h7164; wi = 16'hED38; end
            8'hF5: begin wr = 16'h712B; wi = 16'hEEC6; end
            8'hF6: begin wr = 16'h70F7; wi = 16'hF055; end
            8'hF7: begin wr = 16'h70C9; wi = 16'hF1E4; end
            8'hF8: begin wr = 16'h709F; wi = 16'hF374; end
            8'hF9: begin wr = 16'h807A; wi = 16'hF505; end
            8'hFA: begin wr = 16'h805A; wi = 16'hF696; end
            8'hFB: begin wr = 16'h803F; wi = 16'hF827; end
            8'hFC: begin wr = 16'h8028; wi = 16'hF9B8; end
            8'hFD: begin wr = 16'h8017; wi = 16'hFB4A; end
            8'hFE: begin wr = 16'h800B; wi = 16'hFCDC; end
            8'hFF: begin wr = 16'h8003; wi = 16'hFE6E; end
            default: begin wr = 16'h7FFF; wi = 16'h0000; end
        endcase
    end
endmodule
